package ALU_TYPE is
  type TYPE_OP is (ADD, 
						 ADDC,
						 SUB,
						 SUBC,
						 SUBY,
						 BITAND,
						 BITOR,
						 BITXOR,
						 SL0,
						 SL1,
						 SL_A,
						 SLX,
						 SLC,
						 SR0,
						 SR1,
						 SR_A,
						 SRX,
						 SRC,
						 RR,
						 RL,
						 LOAD,	
						 NOP
						 );

end ALU_TYPE;
                
